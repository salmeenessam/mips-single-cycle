`timescale 1ns / 1ps
module and_gate(
    input A,
    input B,
    output out
    );

assign out = A&B;

endmodule
