`timescale 1ns / 1ps

module and(
    input A,
    input B,
    output out
    );


endmodule
